
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
	    case (Address[9:2])
			0: Instruction <= 32'b00001000000000000000000000010000; // jump to normal入口，第一条jal，然后跳到前面，最后一条jr使得最高位清零
			1: Instruction <= 32'b00001000000000000000000000110000; //jump to Interrupt
			15: Instruction <= 32'b00000011111000000000000000001000;//	jr $ra, $ra中存着17地址
			
			
			16: Instruction <= 32'b000011_00000000000000000000001111;// jal 15
			17: Instruction <= 32'b00111100000011010100000000000000; //gcd代码开始
			18: Instruction <= 32'b10101101101000000000000000001000;
			19: Instruction <= 32'b10101101101000000000000000000000;
			20: Instruction <= 32'b00000000000000000111000000100111;
			21: Instruction <= 32'b10101101101011100000000000000100;
			22: Instruction <= 32'b00100000000011000000000000000011;
			23: Instruction <= 32'b10101101101011000000000000001000;
			24: Instruction <= 32'b00000000000100000100000000101010;
			25: Instruction <= 32'b00000000000100010100100000101010;
			26: Instruction <= 32'b00000001000010010101000000100100;
			27: Instruction <= 32'b00010101010000000000000000000100;
			28: Instruction <= 32'b00000010000000001001000000100000;
			29: Instruction <= 32'b00001000000000000000000000011000;
			30: Instruction <= 32'b00000000000000000000000000000000;
			31: Instruction <= 32'b00000010001000001001100000100000;
			32: Instruction <= 32'b00000010010100110101100000101010;
			33: Instruction <= 32'b00010001011000000000000000000101;
			34: Instruction <= 32'b00000000000000000000000000000000;
			35: Instruction <= 32'b00000010010000000110000000100000;
			36: Instruction <= 32'b00000010011000001001000000100000;
			37: Instruction <= 32'b00000001100000001001100000100000;
			38: Instruction <= 32'b00000010010100111010000000100010;
			39: Instruction <= 32'b00010010100000000000000000000110;
			40: Instruction <= 32'b00000000000000000000000000000000;
			41: Instruction <= 32'b00000010011000001001000000100000;
			42: Instruction <= 32'b00000010100000001001100000100000;
			43: Instruction <= 32'b00001000000000000000000000100000;
			44: Instruction <= 32'b00000000000000000000000000000000;
			45: Instruction <= 32'b10101101101100110000000000011000;
			46: Instruction <= 32'b10101101101100110000000000001100;

			48: Instruction <= 32'b00111100000010000100000000000000;
			49:	Instruction <= 32'b10001101000010010000000000100000;
			50:	Instruction <= 32'b00000000000000000000000000000000;
			51:	Instruction <= 32'b00110001001010100000000000001000;
			52:	Instruction <= 32'b00010001010000000000000000001000;
			53:	Instruction <= 32'b00000000000000000000000000000000;
			54:	Instruction <= 32'b00010010000000000000000000000101;
			55:	Instruction <= 32'b00000000000000000000000000000000;
			56:	Instruction <= 32'b10001101000100010000000000011100;
			57:	Instruction <= 32'b00001000000000000000000000001100;
			58:	Instruction <= 32'b00000000000000000000000000000000;
			59:	Instruction <= 32'b10001101000100000000000000011100;
			60:	Instruction <= 32'b10001101000010010000000000010100;
			61:	Instruction <= 32'b00000000000100010110000100000010;
			62:	Instruction <= 32'b00110001001010100000000100000000;
			63:	Instruction <= 32'b00010001010000000000000000000101;
			64:	Instruction <= 32'b00000000000000000000000000000000;
			65:	Instruction <= 32'b00100000000010110000001000000000;
			66:	Instruction <= 32'b00001000000000000000000000100100;
			67:	Instruction <= 32'b00000000000000000000000000000000;
			68:	Instruction <= 32'b00110001001010100000001000000000;
			69:	Instruction <= 32'b00010001010000000000000000000110;
			70:	Instruction <= 32'b00000000000000000000000000000000;
			71:	Instruction <= 32'b00100000000010110000010000000000;
			72:	Instruction <= 32'b00110010000011000000000000001111;
			73:	Instruction <= 32'b00001000000000000000000000100100;
			74:	Instruction <= 32'b00000000000000000000000000000000;
			75:	Instruction <= 32'b00110001001010100000010000000000;
			76:	Instruction <= 32'b00010001010010010000000000000110;
			77:	Instruction <= 32'b00000000000000000000000000000000;
			78:	Instruction <= 32'b00100000000010110000100000000000;
			79:	Instruction <= 32'b00000000000100000110000100000010;
			80:	Instruction <= 32'b00001000000000000000000000100100;
			81:	Instruction <= 32'b00000000000000000000000000000000;
			82:	Instruction <= 32'b00100000000010110000000100000000;
			83:	Instruction <= 32'b00110010001011000000000000001111;
			84:	Instruction <= 32'b10001101100011010000000000000000;
			85:	Instruction <= 32'b00000000000000000000000000000000;
			86:	Instruction <= 32'b00000001101010110111000000100000;
			87:	Instruction <= 32'b10101101000011100000000000010100;
			88:	Instruction <= 32'b00000011010000000000000000001000;
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
