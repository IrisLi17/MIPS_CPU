`timescale 1ns/1ps

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 64;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin
        ROMDATA[0] <= 32'b00111100000010000100000000000000;
        ROMDATA[1] <= 32'b10001101000010010000000000100000;
        ROMDATA[2] <= 32'b00000000000000000000000000000000;
        ROMDATA[3] <= 32'b00110001001010100000000000001000;
        ROMDATA[4] <= 32'b00010001010000000000000000001000;
        ROMDATA[5] <= 32'b00000000000000000000000000000000;
        ROMDATA[6] <= 32'b00010010000000000000000000000101;
        ROMDATA[7] <= 32'b00000000000000000000000000000000;
        ROMDATA[8] <= 32'b10001101000100010000000000011100;
        ROMDATA[9] <= 32'b00001000000000000000000000001100;
        ROMDATA[10] <= 32'b00000000000000000000000000000000;
        ROMDATA[11] <= 32'b10001101000100000000000000011100;
        ROMDATA[12] <= 32'b10001101000010010000000000010100;
        ROMDATA[13] <= 32'b00000000000100010110000100000010;
        ROMDATA[14] <= 32'b00110001001010100000000100000000;
        ROMDATA[15] <= 32'b00010001010000000000000000000101;
        ROMDATA[16] <= 32'b00000000000000000000000000000000;
        ROMDATA[17] <= 32'b00100000000010110000001000000000;
        ROMDATA[18] <= 32'b00001000000000000000000000100100;
        ROMDATA[19] <= 32'b00000000000000000000000000000000;
        ROMDATA[20] <= 32'b00110001001010100000001000000000;
        ROMDATA[21] <= 32'b00010001010000000000000000000110;
        ROMDATA[22] <= 32'b00000000000000000000000000000000;
        ROMDATA[23] <= 32'b00100000000010110000010000000000;
        ROMDATA[24] <= 32'b00110010000011000000000000001111;
        ROMDATA[25] <= 32'b00001000000000000000000000100100;
        ROMDATA[26] <= 32'b00000000000000000000000000000000;
        ROMDATA[27] <= 32'b00110001001010100000010000000000;
        ROMDATA[28] <= 32'b00010001010010010000000000000110;
        ROMDATA[29] <= 32'b00000000000000000000000000000000;
        ROMDATA[30] <= 32'b00100000000010110000100000000000;
        ROMDATA[31] <= 32'b00000000000100000110000100000010;
        ROMDATA[32] <= 32'b00001000000000000000000000100100;
        ROMDATA[33] <= 32'b00000000000000000000000000000000;
        ROMDATA[34] <= 32'b00100000000010110000000100000000;
        ROMDATA[35] <= 32'b00110010001011000000000000001111;
        ROMDATA[36] <= 32'b10001101100011010000000000000000;
        ROMDATA[37] <= 32'b00000000000000000000000000000000;
        ROMDATA[38] <= 32'b00000001101010110111000000100000;
        ROMDATA[39] <= 32'b10101101000011100000000000010100;
        ROMDATA[40] <= 32'b00000011010000000000000000001000;
	    for (i=41;i<ROM_SIZE;i=i+1) begin
            ROMDATA[i] <= 32'b0;
        end
end
endmodule