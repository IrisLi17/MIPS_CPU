
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
	    case (Address[9:2])
			0: Instruction <= 32'b00001000000000000000000000010000; // jump to normal入口，第�??条jal，然后跳到前面，�??后一条jr使得�??高位清零
			1: Instruction <= 32'b00001000000000000000000001100000; //jump to Interrupt
			2: Instruction <= 32'b00001000000000000000000010100000; // jump to error
			15: Instruction <= 32'b00000011111000000000000000001000;//	jr $ra, $ra中存�??17地址			
			16: Instruction <= 32'b000011_00000000000000000000001111;// jal 15
17: Instruction <= 32'b00111100000011010100000000000000; // ['', ['lui', '$t5', '0x4000']]
18: Instruction <= 32'b10101101101000000000000000001000; // ['', ['sw', '$zero', '8($t5)']]
19: Instruction <= 32'b00111100000011001111111111111111; // ['', ['lui', '$t4', '0xFFFF']]
20: Instruction <= 32'b00100000000011001100000000000000; // ['', ['addi', '$t4', '$zero', '0xFF00']]
21: Instruction <= 32'b10101101101011000000000000000000; // ['', ['sw', '$t4', '0($t5)']]
22: Instruction <= 32'b00000000000000000111000000100111; // ['', ['nor', '$t6', '$zero', '$zero']]
23: Instruction <= 32'b10101101101011100000000000000100; // ['', ['sw', '$t6', '4($t5)']]
24: Instruction <= 32'b00100000000011000000000000000011; // ['', ['addi', '$t4', '$zero', '0x0003']]
25: Instruction <= 32'b10101101101011000000000000001000; // ['', ['sw', '$t4', '8($t5)']]
26: Instruction <= 32'b00000000000101010100000000101010; // ['loop', ['slt', '$t0', '$zero', '$s5']]
27: Instruction <= 32'b00000000000101100100100000101010; // ['', ['slt', '$t1', '$zero', '$s6']]
28: Instruction <= 32'b00000001000010010101000000100100; // ['', ['and', '$t2', '$t0', '$t1']]
29: Instruction <= 32'b00010101010000000000000000000011; // ['', ['bne', '$t2', '$zero', 'target']]
30: Instruction <= 32'b00000010101000001001000000100000; // ['', ['add', '$s2', '$s5', '$zero']]
31: Instruction <= 32'b00001000000000000000000000011010; // ['', ['j', 'loop']]
32: Instruction <= 32'b00000000000000000000000000000000; // ['', ['sll', '$zero', '$zero', '0']]
33: Instruction <= 32'b00000010110000001001100000100000; // ['target', ['add', '$s3', '$s6', '$zero']]
34: Instruction <= 32'b00000010010100110101100000101010; // ['compare', ['slt', '$t3', '$s2', '$s3']]
35: Instruction <= 32'b00010001011000000000000000000100; // ['', ['beq', '$t3', '$zero', 's2greater']]
36: Instruction <= 32'b00000000000000000000000000000000; // ['', ['sll', '$zero', '$zero', '0']]
37: Instruction <= 32'b00000010010000000110000000100000; // ['', ['add', '$t4', '$s2', '$zero']]
38: Instruction <= 32'b00000010011000001001000000100000; // ['', ['add', '$s2', '$s3', '$zero']]
39: Instruction <= 32'b00000001100000001001100000100000; // ['', ['add', '$s3', '$t4', '$zero']]
40: Instruction <= 32'b00000010010100111010000000100010; // ['s2greater', ['sub', '$s4', '$s2', '$s3']]
41: Instruction <= 32'b00010010100000000000000000000101; // ['', ['beq', '$s4', '$zero', 'finish']]
42: Instruction <= 32'b00000000000000000000000000000000; // ['', ['sll', '$zero', '$zero', '0']]
43: Instruction <= 32'b00000010011000001001000000100000; // ['', ['add', '$s2', '$s3', '$zero']]
44: Instruction <= 32'b00000010100000001001100000100000; // ['', ['add', '$s3', '$s4', '$zero']]
45: Instruction <= 32'b00001000000000000000000000100010; // ['', ['j', 'compare']]
46: Instruction <= 32'b00000000000000000000000000000000; // ['', ['sll', '$zero', '$zero', '0']]
47: Instruction <= 32'b00111100000011010100000000000000; // ['finish', ['lui', '$t5', '0x4000']]
48: Instruction <= 32'b10101101101100110000000000011000; // ['', ['sw', '$s3', '24($t5)']]
49: Instruction <= 32'b10101101101100110000000000001100; // ['', ['sw', '$s3', '12($t5)']]
50: Instruction <= 32'b00000000000000001010100000100000; // ['', ['add', '$s5', '$zero', '$zero']]
51: Instruction <= 32'b00000000000000001011000000100000; // ['', ['add', '$s6', '$zero', '$zero']]
52: Instruction <= 32'b00001000000000000000000000110101; // ['', ['j', 'Exit']]
53: Instruction <= 32'b00111100000010000100000000000000; // ['Exit', ['lui', '$t0', '0x4000']]
54: Instruction <= 32'b10001101000010010000000000100000; // ['', ['lw', '$t1', '32($t0)']]
55: Instruction <= 32'b00100000000010100000000000001000; // ['', ['addi', '$t2', '$zero', '8']]
56: Instruction <= 32'b00000001001010100100100000100100; // ['', ['and', '$t1', '$t1', '$t2']]
57: Instruction <= 32'b00010101001000001111111111100000; // ['', ['bne', '$t1', '$zero', 'loop']]
58: Instruction <= 32'b00001000000000000000000000110101; // ['', ['j', 'Exit']]


96: Instruction <= 32'b00100011101111011111111111100100; // ['', ['addi', '$sp', '$sp', '-28']]
97: Instruction <= 32'b10101111101011100000000000011000; // ['', ['sw', '$t6', '24($sp)']]
98: Instruction <= 32'b10101111101011010000000000010100; // ['', ['sw', '$t5', '20($sp)']]
99: Instruction <= 32'b10101111101011000000000000010000; // ['', ['sw', '$t4', '16($sp)']]
100: Instruction <= 32'b10101111101010110000000000001100; // ['', ['sw', '$t3', '12($sp)']]
101: Instruction <= 32'b10101111101010100000000000001000; // ['', ['sw', '$t2', '8($sp)']]
102: Instruction <= 32'b10101111101010010000000000000100; // ['', ['sw', '$t1', '4($sp)']]
103: Instruction <= 32'b10101111101010000000000000000000; // ['', ['sw', '$t0', '0($sp)']]
104: Instruction <= 32'b00111100000010000100000000000000; // ['', ['lui', '$t0', '0x4000']]
105: Instruction <= 32'b10001101000010010000000000001000; // ['', ['lw', '$t1', '8($t0)']]
106: Instruction <= 32'b00100000000010101111111111111001; // ['', ['addi', '$t2', '$zero', '0xFFF9']]
107: Instruction <= 32'b00000001001010100100100000100100; // ['', ['and', '$t1', '$t1', '$t2']]
108: Instruction <= 32'b10101101000010010000000000001000; // ['', ['sw', '$t1', '8($t0)']]
109: Instruction <= 32'b10001101000010010000000000100000; // ['', ['lw', '$t1', '32($t0)']]
110: Instruction <= 32'b00110001001010100000000000001000; // ['', ['andi', '$t2', '$t1', '0x0008']]
111: Instruction <= 32'b00010001010000000000000000000111; // ['', ['beq', '$t2', '$zero', 'noload']]
112: Instruction <= 32'b00010010101000000000000000000100; // ['', ['beq', '$s5', '$zero', 'loads0']]
113: Instruction <= 32'b00010110110000000000000000000101; // ['', ['bne', '$s6', '$zero', 'noload']]
114: Instruction <= 32'b10001101000100010000000000011100; // ['', ['lw', '$s1', '28($t0)']]
115: Instruction <= 32'b00100010001101100000000000000000; // ['', ['addi', '$s6', '$s1', '0']]
116: Instruction <= 32'b00001000000000000000000001110111; // ['', ['j', 'noload']]
117: Instruction <= 32'b10001101000100000000000000011100; // ['loads0', ['lw', '$s0', '28($t0)']]
118: Instruction <= 32'b00100010000101010000000000000000; // ['', ['addi', '$s5', '$s0', '0']]
119: Instruction <= 32'b10001101000010010000000000010100; // ['noload', ['lw', '$t1', '20($t0)']]
120: Instruction <= 32'b00000000000100010110000100000010; // ['', ['srl', '$t4', '$s1', '4']]
121: Instruction <= 32'b00110001001010100000000100000000; // ['', ['andi', '$t2', '$t1', '0x0100']]
122: Instruction <= 32'b00010001010000000000000000000010; // ['', ['beq', '$t2', '$zero', 'target1']]
123: Instruction <= 32'b00100000000010110000001000000000; // ['', ['addi', '$t3', '$zero', '0x0200']]
124: Instruction <= 32'b00001000000000000000000010001001; // ['', ['j', 'finish']]
125: Instruction <= 32'b00110001001010100000001000000000; // ['target1', ['andi', '$t2', '$t1', '0x0200']]
126: Instruction <= 32'b00010001010000000000000000000011; // ['', ['beq', '$t2', '$zero', 'target2']]
127: Instruction <= 32'b00100000000010110000010000000000; // ['', ['addi', '$t3', '$zero', '0x0400']]
128: Instruction <= 32'b00110010000011000000000000001111; // ['', ['andi', '$t4', '$s0', '0x000F']]
129: Instruction <= 32'b00001000000000000000000010001001; // ['', ['j', 'finish']]
130: Instruction <= 32'b00110001001010100000010000000000; // ['target2', ['andi', '$t2', '$t1', '0x0400']]
131: Instruction <= 32'b00010001010000000000000000000011; // ['', ['beq', '$t2', '$zero', 'target3']]
132: Instruction <= 32'b00100000000010110000100000000000; // ['', ['addi', '$t3', '$zero', '0x0800']]
133: Instruction <= 32'b00000000000100000110000100000010; // ['', ['srl', '$t4', '$s0', '4']]
134: Instruction <= 32'b00001000000000000000000010001001; // ['', ['j', 'finish']]
135: Instruction <= 32'b00100000000010110000000100000000; // ['target3', ['addi', '$t3', '$zero', '0x0100']]
136: Instruction <= 32'b00110010001011000000000000001111; // ['', ['andi', '$t4', '$s1', '0x000F']]
137: Instruction <= 32'b00000000000011000110000010000000; // ['finish', ['sll', '$t4', '$t4', '2']]
138: Instruction <= 32'b10001101100011010000000000000000; // ['', ['lw', '$t5', '0($t4)']]
139: Instruction <= 32'b00000001101010110111000000100000; // ['', ['add', '$t6', '$t5', '$t3']]
140: Instruction <= 32'b10101101000011100000000000010100; // ['', ['sw', '$t6', '20($t0)']]
141: Instruction <= 32'b10001101000010010000000000001000; // ['', ['lw', '$t1', '8($t0)']]
142: Instruction <= 32'b00100000000010100000000000000010; // ['', ['addi', '$t2', '$zero', '0x0002']]
143: Instruction <= 32'b00000001001010100101100000100101; // ['', ['or', '$t3', '$t1', '$t2']]
144: Instruction <= 32'b10101101000010110000000000001000; // ['', ['sw', '$t3', '8($t0)']]
145: Instruction <= 32'b10001111101010000000000000000000; // ['', ['lw', '$t0', '0($sp)']]
146: Instruction <= 32'b10001111101010010000000000000100; // ['', ['lw', '$t1', '4($sp)']]
147: Instruction <= 32'b10001111101010100000000000001000; // ['', ['lw', '$t2', '8($sp)']]
148: Instruction <= 32'b10001111101010110000000000001100; // ['', ['lw', '$t3', '12($sp)']]
149: Instruction <= 32'b10001111101011000000000000010000; // ['', ['lw', '$t4', '16($sp)']]
150: Instruction <= 32'b10001111101011010000000000010100; // ['', ['lw', '$t5', '20($sp)']]
151: Instruction <= 32'b10001111101011100000000000011000; // ['', ['lw', '$t6', '24($sp)']]
152: Instruction <= 32'b00100011101111010000000000011100; // ['', ['addi', '$sp', '$sp', '28']]
153: Instruction <= 32'b00000011010000000000000000001000; // ['', ['jr', '$k0']]

160: Instruction <= 32'b00000000000000000000000000000000; // ['error', ['nop']]
161: Instruction <= 32'b00001000000000000000000010100000; // ['', ['j', 'error']] 
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
