
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
	    case (Address[9:2])
			0: Instruction <= 32'b00001000000000000000000000010000; // jump to normal入口，第一条jal，然后跳到前面，最后一条jr使得最高位清零
			1: Instruction <= 32'b00001000000000000000000001100000; //jump to Interrupt
			15: Instruction <= 32'b00000011111000000000000000001000;//	jr $ra, $ra中存着17地址
			
			
			16: Instruction <= 32'b000011_00000000000000000000001111;// jal 15
17: Instruction <= 32'b00111100000011010100000000000000; // gcd begin
18: Instruction <= 32'b10101101101000000000000000001000;
19: Instruction <= 32'b00111100000011001111111111111111;
20: Instruction <= 32'b00100000000011001111000000000000;
21: Instruction <= 32'b10101101101011000000000000000000;
22: Instruction <= 32'b00000000000000000111000000100111;
23: Instruction <= 32'b10101101101011100000000000000100;
24: Instruction <= 32'b00100000000011000000000000000011;
25: Instruction <= 32'b10101101101011000000000000001000;
26: Instruction <= 32'b00000000000100000100000000101010;
27: Instruction <= 32'b00000000000100010100100000101010;
28: Instruction <= 32'b00000001000010010101000000100100;
29: Instruction <= 32'b00010101010000000000000000000100;
30: Instruction <= 32'b00000010000000001001000000100000;
31: Instruction <= 32'b00001000000000000000000000011010;
32: Instruction <= 32'b00000000000000000000000000000000;
33: Instruction <= 32'b00000010001000001001100000100000;
34: Instruction <= 32'b00000010010100110101100000101010;
35: Instruction <= 32'b00010001011000000000000000000100;
36: Instruction <= 32'b00000000000000000000000000000000;
37: Instruction <= 32'b00000010010000000110000000100000;
38: Instruction <= 32'b00000010011000001001000000100000;
39: Instruction <= 32'b00000001100000001001100000100000;
40: Instruction <= 32'b00000010010100111010000000100010;
41: Instruction <= 32'b00010010100000000000000000000101;
42: Instruction <= 32'b00000000000000000000000000000000;
43: Instruction <= 32'b00000010011000001001000000100000;
44: Instruction <= 32'b00000010100000001001100000100000;
45: Instruction <= 32'b00001000000000000000000000100010;
46: Instruction <= 32'b00000000000000000000000000000000;
47: Instruction <= 32'b10101101101100110000000000011000;
48: Instruction <= 32'b10101101101100110000000000001100;


96: Instruction <= 32'b00100011101111010000000000011100;
97: Instruction <= 32'b10101111101011100000000000011000;
98: Instruction <= 32'b10101111101011010000000000010100;
99: Instruction <= 32'b10101111101011000000000000010000;
100: Instruction <= 32'b10101111101010110000000000001100;
101: Instruction <= 32'b10101111101010100000000000001000;
102: Instruction <= 32'b10101111101010010000000000000100;
103: Instruction <= 32'b10101111101010000000000000000000;
104: Instruction <= 32'b00111100000010000100000000000000;
105: Instruction <= 32'b10001101000010010000000000001000;
106: Instruction <= 32'b00100000000010101111111111111001;
107: Instruction <= 32'b00000001001010100100100000100100;
108: Instruction <= 32'b10101101000010010000000000001000;
109: Instruction <= 32'b10001101000010010000000000100000;
110: Instruction <= 32'b00110001001010100000000000001000;
111: Instruction <= 32'b00010001010000000000000000000100;
112: Instruction <= 32'b00010010000000000000000000000010;
113: Instruction <= 32'b10001101000100010000000000011100;
114: Instruction <= 32'b00001000000000000000000001110100;
115: Instruction <= 32'b10001101000100000000000000011100;
116: Instruction <= 32'b10001101000010010000000000010100;
117: Instruction <= 32'b00000000000100010110000100000010;
118: Instruction <= 32'b00110001001010100000000100000000;
119: Instruction <= 32'b00010001010000000000000000000010;
120: Instruction <= 32'b00100000000010110000001000000000;
121: Instruction <= 32'b00001000000000000000000010000110;
122: Instruction <= 32'b00110001001010100000001000000000;
123: Instruction <= 32'b00010001010000000000000000000011;
124: Instruction <= 32'b00100000000010110000010000000000;
125: Instruction <= 32'b00110010000011000000000000001111;
126: Instruction <= 32'b00001000000000000000000010000110;
127: Instruction <= 32'b00110001001010100000010000000000;
128: Instruction <= 32'b00010001010010010000000000000011;
129: Instruction <= 32'b00100000000010110000100000000000;
130: Instruction <= 32'b00000000000100000110000100000010;
131: Instruction <= 32'b00001000000000000000000010000110;
132: Instruction <= 32'b00100000000010110000000100000000;
133: Instruction <= 32'b00110010001011000000000000001111;
134: Instruction <= 32'b10001101100011010000000000000000;
135: Instruction <= 32'b00000001101010110111000000100000;
136: Instruction <= 32'b10101101000011100000000000010100;
137: Instruction <= 32'b10001101000010010000000000001000;
138: Instruction <= 32'b00100000000010100000000000000010;
139: Instruction <= 32'b00000001001010100101100000100101;
140: Instruction <= 32'b10101101000010110000000000001000;
141: Instruction <= 32'b10001111101010000000000000000000;
142: Instruction <= 32'b10001101001010010000000000000100;
143: Instruction <= 32'b10001111101010100000000000001000;
144: Instruction <= 32'b10001111101010110000000000001100;
145: Instruction <= 32'b10001111101011000000000000010000;
146: Instruction <= 32'b10001111101011010000000000010100;
147: Instruction <= 32'b10001111101011100000000000011000;
148: Instruction <= 32'b00100011101111010000000000011100;
149: Instruction <= 32'b00000011010000000000000000001000;

			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
